// platform.v

// Generated using ACDS version 19.1 670

`timescale 1 ps / 1 ps
module platform (
		input  wire        clk_clk,          //        clk.clk
		output wire [9:0]  ledr_export,      //       ledr.export
		input  wire        reset_reset,      //      reset.reset
		output wire        sdram_clk_clk,    //  sdram_clk.clk
		output wire [12:0] sdram_wire_addr,  // sdram_wire.addr
		output wire [1:0]  sdram_wire_ba,    //           .ba
		output wire        sdram_wire_cas_n, //           .cas_n
		output wire        sdram_wire_cke,   //           .cke
		output wire        sdram_wire_cs_n,  //           .cs_n
		inout  wire [15:0] sdram_wire_dq,    //           .dq
		output wire [1:0]  sdram_wire_dqm,   //           .dqm
		output wire        sdram_wire_ras_n, //           .ras_n
		output wire        sdram_wire_we_n,  //           .we_n
		input  wire [9:0]  sw_export         //         sw.export
	);

	wire  [31:0] riscv_simple_sv_0_text_master_readdata;         // Instruction_Cache_0:core_instruction -> riscv_simple_sv_0:inst_data
	wire         riscv_simple_sv_0_text_master_waitrequest;      // Instruction_Cache_0:core_waitrequest -> riscv_simple_sv_0:inst_wait_req
	wire  [31:0] riscv_simple_sv_0_text_master_address;          // riscv_simple_sv_0:pc -> Instruction_Cache_0:core_inst_address
	wire         riscv_simple_sv_0_text_master_read;             // riscv_simple_sv_0:inst_read_enable -> Instruction_Cache_0:core_read
	wire         riscv_simple_sv_0_text_master_readdatavalid;    // Instruction_Cache_0:core_inst_valid -> riscv_simple_sv_0:inst_valid
	wire         sys_sdram_pll_sys_clk_clk;                      // sys_sdram_pll:sys_clk_clk -> [Instruction_Cache_0:clock, jtag_master:clk_clk, ledr:clk, mm_interconnect_0:sys_sdram_pll_sys_clk_clk, riscv_data:clk, riscv_sdram:clk, riscv_simple_sv_0:clock, riscv_text:clk, rst_controller:clk, rst_controller_001:clk, sw:clk]
	wire         sys_sdram_pll_reset_source_reset;               // sys_sdram_pll:reset_source_reset -> [jtag_master:clk_reset_reset, rst_controller:reset_in0, rst_controller_001:reset_in1]
	wire  [31:0] riscv_simple_sv_0_data_master_readdata;         // mm_interconnect_0:riscv_simple_sv_0_data_master_readdata -> riscv_simple_sv_0:bus_read_data
	wire         riscv_simple_sv_0_data_master_waitrequest;      // mm_interconnect_0:riscv_simple_sv_0_data_master_waitrequest -> riscv_simple_sv_0:bus_wait_req
	wire  [31:0] riscv_simple_sv_0_data_master_address;          // riscv_simple_sv_0:bus_address -> mm_interconnect_0:riscv_simple_sv_0_data_master_address
	wire   [3:0] riscv_simple_sv_0_data_master_byteenable;       // riscv_simple_sv_0:bus_byte_enable -> mm_interconnect_0:riscv_simple_sv_0_data_master_byteenable
	wire         riscv_simple_sv_0_data_master_read;             // riscv_simple_sv_0:bus_read_enable -> mm_interconnect_0:riscv_simple_sv_0_data_master_read
	wire         riscv_simple_sv_0_data_master_readdatavalid;    // mm_interconnect_0:riscv_simple_sv_0_data_master_readdatavalid -> riscv_simple_sv_0:bus_valid
	wire  [31:0] riscv_simple_sv_0_data_master_writedata;        // riscv_simple_sv_0:bus_write_data -> mm_interconnect_0:riscv_simple_sv_0_data_master_writedata
	wire         riscv_simple_sv_0_data_master_write;            // riscv_simple_sv_0:bus_write_enable -> mm_interconnect_0:riscv_simple_sv_0_data_master_write
	wire  [31:0] jtag_master_master_readdata;                    // mm_interconnect_0:jtag_master_master_readdata -> jtag_master:master_readdata
	wire         jtag_master_master_waitrequest;                 // mm_interconnect_0:jtag_master_master_waitrequest -> jtag_master:master_waitrequest
	wire  [31:0] jtag_master_master_address;                     // jtag_master:master_address -> mm_interconnect_0:jtag_master_master_address
	wire         jtag_master_master_read;                        // jtag_master:master_read -> mm_interconnect_0:jtag_master_master_read
	wire   [3:0] jtag_master_master_byteenable;                  // jtag_master:master_byteenable -> mm_interconnect_0:jtag_master_master_byteenable
	wire         jtag_master_master_readdatavalid;               // mm_interconnect_0:jtag_master_master_readdatavalid -> jtag_master:master_readdatavalid
	wire         jtag_master_master_write;                       // jtag_master:master_write -> mm_interconnect_0:jtag_master_master_write
	wire  [31:0] jtag_master_master_writedata;                   // jtag_master:master_writedata -> mm_interconnect_0:jtag_master_master_writedata
	wire  [63:0] instruction_cache_0_memory_readdata;            // mm_interconnect_0:Instruction_Cache_0_memory_readdata -> Instruction_Cache_0:memory_readdata
	wire         instruction_cache_0_memory_waitrequest;         // mm_interconnect_0:Instruction_Cache_0_memory_waitrequest -> Instruction_Cache_0:memory_waitrequest
	wire  [31:0] instruction_cache_0_memory_address;             // Instruction_Cache_0:memory_address -> mm_interconnect_0:Instruction_Cache_0_memory_address
	wire         instruction_cache_0_memory_read;                // Instruction_Cache_0:memory_read -> mm_interconnect_0:Instruction_Cache_0_memory_read
	wire         instruction_cache_0_memory_readdatavalid;       // mm_interconnect_0:Instruction_Cache_0_memory_readdatavalid -> Instruction_Cache_0:memory_readdatavalid
	wire   [3:0] instruction_cache_0_memory_burstcount;          // Instruction_Cache_0:memory_burstcount -> mm_interconnect_0:Instruction_Cache_0_memory_burstcount
	wire         mm_interconnect_0_riscv_sdram_s1_chipselect;    // mm_interconnect_0:riscv_sdram_s1_chipselect -> riscv_sdram:az_cs
	wire  [15:0] mm_interconnect_0_riscv_sdram_s1_readdata;      // riscv_sdram:za_data -> mm_interconnect_0:riscv_sdram_s1_readdata
	wire         mm_interconnect_0_riscv_sdram_s1_waitrequest;   // riscv_sdram:za_waitrequest -> mm_interconnect_0:riscv_sdram_s1_waitrequest
	wire  [24:0] mm_interconnect_0_riscv_sdram_s1_address;       // mm_interconnect_0:riscv_sdram_s1_address -> riscv_sdram:az_addr
	wire         mm_interconnect_0_riscv_sdram_s1_read;          // mm_interconnect_0:riscv_sdram_s1_read -> riscv_sdram:az_rd_n
	wire   [1:0] mm_interconnect_0_riscv_sdram_s1_byteenable;    // mm_interconnect_0:riscv_sdram_s1_byteenable -> riscv_sdram:az_be_n
	wire         mm_interconnect_0_riscv_sdram_s1_readdatavalid; // riscv_sdram:za_valid -> mm_interconnect_0:riscv_sdram_s1_readdatavalid
	wire         mm_interconnect_0_riscv_sdram_s1_write;         // mm_interconnect_0:riscv_sdram_s1_write -> riscv_sdram:az_wr_n
	wire  [15:0] mm_interconnect_0_riscv_sdram_s1_writedata;     // mm_interconnect_0:riscv_sdram_s1_writedata -> riscv_sdram:az_data
	wire         mm_interconnect_0_ledr_s1_chipselect;           // mm_interconnect_0:ledr_s1_chipselect -> ledr:chipselect
	wire  [31:0] mm_interconnect_0_ledr_s1_readdata;             // ledr:readdata -> mm_interconnect_0:ledr_s1_readdata
	wire   [1:0] mm_interconnect_0_ledr_s1_address;              // mm_interconnect_0:ledr_s1_address -> ledr:address
	wire         mm_interconnect_0_ledr_s1_write;                // mm_interconnect_0:ledr_s1_write -> ledr:write_n
	wire  [31:0] mm_interconnect_0_ledr_s1_writedata;            // mm_interconnect_0:ledr_s1_writedata -> ledr:writedata
	wire  [31:0] mm_interconnect_0_sw_s1_readdata;               // sw:readdata -> mm_interconnect_0:sw_s1_readdata
	wire   [1:0] mm_interconnect_0_sw_s1_address;                // mm_interconnect_0:sw_s1_address -> sw:address
	wire         mm_interconnect_0_riscv_text_s1_chipselect;     // mm_interconnect_0:riscv_text_s1_chipselect -> riscv_text:chipselect
	wire  [31:0] mm_interconnect_0_riscv_text_s1_readdata;       // riscv_text:readdata -> mm_interconnect_0:riscv_text_s1_readdata
	wire  [13:0] mm_interconnect_0_riscv_text_s1_address;        // mm_interconnect_0:riscv_text_s1_address -> riscv_text:address
	wire   [3:0] mm_interconnect_0_riscv_text_s1_byteenable;     // mm_interconnect_0:riscv_text_s1_byteenable -> riscv_text:byteenable
	wire         mm_interconnect_0_riscv_text_s1_write;          // mm_interconnect_0:riscv_text_s1_write -> riscv_text:write
	wire  [31:0] mm_interconnect_0_riscv_text_s1_writedata;      // mm_interconnect_0:riscv_text_s1_writedata -> riscv_text:writedata
	wire         mm_interconnect_0_riscv_text_s1_clken;          // mm_interconnect_0:riscv_text_s1_clken -> riscv_text:clken
	wire         mm_interconnect_0_riscv_data_s1_chipselect;     // mm_interconnect_0:riscv_data_s1_chipselect -> riscv_data:chipselect
	wire  [31:0] mm_interconnect_0_riscv_data_s1_readdata;       // riscv_data:readdata -> mm_interconnect_0:riscv_data_s1_readdata
	wire  [14:0] mm_interconnect_0_riscv_data_s1_address;        // mm_interconnect_0:riscv_data_s1_address -> riscv_data:address
	wire   [3:0] mm_interconnect_0_riscv_data_s1_byteenable;     // mm_interconnect_0:riscv_data_s1_byteenable -> riscv_data:byteenable
	wire         mm_interconnect_0_riscv_data_s1_write;          // mm_interconnect_0:riscv_data_s1_write -> riscv_data:write
	wire  [31:0] mm_interconnect_0_riscv_data_s1_writedata;      // mm_interconnect_0:riscv_data_s1_writedata -> riscv_data:writedata
	wire         mm_interconnect_0_riscv_data_s1_clken;          // mm_interconnect_0:riscv_data_s1_clken -> riscv_data:clken
	wire         rst_controller_reset_out_reset;                 // rst_controller:reset_out -> [Instruction_Cache_0:reset, mm_interconnect_0:Instruction_Cache_0_reset_reset_bridge_in_reset_reset, mm_interconnect_0:jtag_master_clk_reset_reset_bridge_in_reset_reset, sw:reset_n]
	wire         rst_controller_001_reset_out_reset;             // rst_controller_001:reset_out -> [ledr:reset_n, mm_interconnect_0:riscv_simple_sv_0_reset_reset_bridge_in_reset_reset, riscv_data:reset, riscv_sdram:reset_n, riscv_simple_sv_0:reset, riscv_text:reset, rst_translator:in_reset]
	wire         rst_controller_001_reset_out_reset_req;         // rst_controller_001:reset_req -> [riscv_data:reset_req, riscv_text:reset_req, rst_translator:reset_req_in]
	wire         jtag_master_master_reset_reset;                 // jtag_master:master_reset_reset -> rst_controller_001:reset_in0

	instruction_cache #(
		.number_of_sets        (4),
		.bits_for_index        (6),
		.bits_for_offset       (6),
		.log_of_number_of_sets (2)
	) instruction_cache_0 (
		.reset                (rst_controller_reset_out_reset),              //  reset.reset
		.core_waitrequest     (riscv_simple_sv_0_text_master_waitrequest),   //   core.waitrequest
		.core_read            (riscv_simple_sv_0_text_master_read),          //       .read
		.core_inst_address    (riscv_simple_sv_0_text_master_address),       //       .address
		.core_instruction     (riscv_simple_sv_0_text_master_readdata),      //       .readdata
		.core_inst_valid      (riscv_simple_sv_0_text_master_readdatavalid), //       .readdatavalid
		.clock                (sys_sdram_pll_sys_clk_clk),                   //  clock.clk
		.memory_address       (instruction_cache_0_memory_address),          // memory.address
		.memory_read          (instruction_cache_0_memory_read),             //       .read
		.memory_readdata      (instruction_cache_0_memory_readdata),         //       .readdata
		.memory_waitrequest   (instruction_cache_0_memory_waitrequest),      //       .waitrequest
		.memory_burstcount    (instruction_cache_0_memory_burstcount),       //       .burstcount
		.memory_readdatavalid (instruction_cache_0_memory_readdatavalid)     //       .readdatavalid
	);

	platform_jtag_master #(
		.USE_PLI     (0),
		.PLI_PORT    (50000),
		.FIFO_DEPTHS (2)
	) jtag_master (
		.clk_clk              (sys_sdram_pll_sys_clk_clk),        //          clk.clk
		.clk_reset_reset      (sys_sdram_pll_reset_source_reset), //    clk_reset.reset
		.master_address       (jtag_master_master_address),       //       master.address
		.master_readdata      (jtag_master_master_readdata),      //             .readdata
		.master_read          (jtag_master_master_read),          //             .read
		.master_write         (jtag_master_master_write),         //             .write
		.master_writedata     (jtag_master_master_writedata),     //             .writedata
		.master_waitrequest   (jtag_master_master_waitrequest),   //             .waitrequest
		.master_readdatavalid (jtag_master_master_readdatavalid), //             .readdatavalid
		.master_byteenable    (jtag_master_master_byteenable),    //             .byteenable
		.master_reset_reset   (jtag_master_master_reset_reset)    // master_reset.reset
	);

	platform_ledr ledr (
		.clk        (sys_sdram_pll_sys_clk_clk),            //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),  //               reset.reset_n
		.address    (mm_interconnect_0_ledr_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_ledr_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_ledr_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_ledr_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_ledr_s1_readdata),   //                    .readdata
		.out_port   (ledr_export)                           // external_connection.export
	);

	platform_riscv_data riscv_data (
		.clk        (sys_sdram_pll_sys_clk_clk),                  //   clk1.clk
		.address    (mm_interconnect_0_riscv_data_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_riscv_data_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_riscv_data_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_riscv_data_s1_write),      //       .write
		.readdata   (mm_interconnect_0_riscv_data_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_riscv_data_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_riscv_data_s1_byteenable), //       .byteenable
		.reset      (rst_controller_001_reset_out_reset),         // reset1.reset
		.reset_req  (rst_controller_001_reset_out_reset_req),     //       .reset_req
		.freeze     (1'b0)                                        // (terminated)
	);

	platform_riscv_sdram riscv_sdram (
		.clk            (sys_sdram_pll_sys_clk_clk),                      //   clk.clk
		.reset_n        (~rst_controller_001_reset_out_reset),            // reset.reset_n
		.az_addr        (mm_interconnect_0_riscv_sdram_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_riscv_sdram_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_riscv_sdram_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_riscv_sdram_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_riscv_sdram_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_riscv_sdram_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_riscv_sdram_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_riscv_sdram_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_riscv_sdram_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_wire_addr),                                //  wire.export
		.zs_ba          (sdram_wire_ba),                                  //      .export
		.zs_cas_n       (sdram_wire_cas_n),                               //      .export
		.zs_cke         (sdram_wire_cke),                                 //      .export
		.zs_cs_n        (sdram_wire_cs_n),                                //      .export
		.zs_dq          (sdram_wire_dq),                                  //      .export
		.zs_dqm         (sdram_wire_dqm),                                 //      .export
		.zs_ras_n       (sdram_wire_ras_n),                               //      .export
		.zs_we_n        (sdram_wire_we_n)                                 //      .export
	);

	riscv_core riscv_simple_sv_0 (
		.reset            (rst_controller_001_reset_out_reset),          //       reset.reset
		.clock            (sys_sdram_pll_sys_clk_clk),                   //       clock.clk
		.pc               (riscv_simple_sv_0_text_master_address),       // text_master.address
		.inst_data        (riscv_simple_sv_0_text_master_readdata),      //            .readdata
		.inst_valid       (riscv_simple_sv_0_text_master_readdatavalid), //            .readdatavalid
		.inst_wait_req    (riscv_simple_sv_0_text_master_waitrequest),   //            .waitrequest
		.inst_read_enable (riscv_simple_sv_0_text_master_read),          //            .read
		.bus_address      (riscv_simple_sv_0_data_master_address),       // data_master.address
		.bus_read_data    (riscv_simple_sv_0_data_master_readdata),      //            .readdata
		.bus_write_data   (riscv_simple_sv_0_data_master_writedata),     //            .writedata
		.bus_byte_enable  (riscv_simple_sv_0_data_master_byteenable),    //            .byteenable
		.bus_read_enable  (riscv_simple_sv_0_data_master_read),          //            .read
		.bus_write_enable (riscv_simple_sv_0_data_master_write),         //            .write
		.bus_wait_req     (riscv_simple_sv_0_data_master_waitrequest),   //            .waitrequest
		.bus_valid        (riscv_simple_sv_0_data_master_readdatavalid)  //            .readdatavalid
	);

	platform_riscv_text riscv_text (
		.clk        (sys_sdram_pll_sys_clk_clk),                  //   clk1.clk
		.address    (mm_interconnect_0_riscv_text_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_riscv_text_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_riscv_text_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_riscv_text_s1_write),      //       .write
		.readdata   (mm_interconnect_0_riscv_text_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_riscv_text_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_riscv_text_s1_byteenable), //       .byteenable
		.reset      (rst_controller_001_reset_out_reset),         // reset1.reset
		.reset_req  (rst_controller_001_reset_out_reset_req),     //       .reset_req
		.freeze     (1'b0)                                        // (terminated)
	);

	platform_sw sw (
		.clk      (sys_sdram_pll_sys_clk_clk),        //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),  //               reset.reset_n
		.address  (mm_interconnect_0_sw_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_sw_s1_readdata), //                    .readdata
		.in_port  (sw_export)                         // external_connection.export
	);

	platform_sys_sdram_pll sys_sdram_pll (
		.ref_clk_clk        (clk_clk),                          //      ref_clk.clk
		.ref_reset_reset    (reset_reset),                      //    ref_reset.reset
		.sys_clk_clk        (sys_sdram_pll_sys_clk_clk),        //      sys_clk.clk
		.sdram_clk_clk      (sdram_clk_clk),                    //    sdram_clk.clk
		.reset_source_reset (sys_sdram_pll_reset_source_reset)  // reset_source.reset
	);

	platform_mm_interconnect_0 mm_interconnect_0 (
		.sys_sdram_pll_sys_clk_clk                             (sys_sdram_pll_sys_clk_clk),                      //                           sys_sdram_pll_sys_clk.clk
		.Instruction_Cache_0_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                 // Instruction_Cache_0_reset_reset_bridge_in_reset.reset
		.jtag_master_clk_reset_reset_bridge_in_reset_reset     (rst_controller_reset_out_reset),                 //     jtag_master_clk_reset_reset_bridge_in_reset.reset
		.riscv_simple_sv_0_reset_reset_bridge_in_reset_reset   (rst_controller_001_reset_out_reset),             //   riscv_simple_sv_0_reset_reset_bridge_in_reset.reset
		.Instruction_Cache_0_memory_address                    (instruction_cache_0_memory_address),             //                      Instruction_Cache_0_memory.address
		.Instruction_Cache_0_memory_waitrequest                (instruction_cache_0_memory_waitrequest),         //                                                .waitrequest
		.Instruction_Cache_0_memory_burstcount                 (instruction_cache_0_memory_burstcount),          //                                                .burstcount
		.Instruction_Cache_0_memory_read                       (instruction_cache_0_memory_read),                //                                                .read
		.Instruction_Cache_0_memory_readdata                   (instruction_cache_0_memory_readdata),            //                                                .readdata
		.Instruction_Cache_0_memory_readdatavalid              (instruction_cache_0_memory_readdatavalid),       //                                                .readdatavalid
		.jtag_master_master_address                            (jtag_master_master_address),                     //                              jtag_master_master.address
		.jtag_master_master_waitrequest                        (jtag_master_master_waitrequest),                 //                                                .waitrequest
		.jtag_master_master_byteenable                         (jtag_master_master_byteenable),                  //                                                .byteenable
		.jtag_master_master_read                               (jtag_master_master_read),                        //                                                .read
		.jtag_master_master_readdata                           (jtag_master_master_readdata),                    //                                                .readdata
		.jtag_master_master_readdatavalid                      (jtag_master_master_readdatavalid),               //                                                .readdatavalid
		.jtag_master_master_write                              (jtag_master_master_write),                       //                                                .write
		.jtag_master_master_writedata                          (jtag_master_master_writedata),                   //                                                .writedata
		.riscv_simple_sv_0_data_master_address                 (riscv_simple_sv_0_data_master_address),          //                   riscv_simple_sv_0_data_master.address
		.riscv_simple_sv_0_data_master_waitrequest             (riscv_simple_sv_0_data_master_waitrequest),      //                                                .waitrequest
		.riscv_simple_sv_0_data_master_byteenable              (riscv_simple_sv_0_data_master_byteenable),       //                                                .byteenable
		.riscv_simple_sv_0_data_master_read                    (riscv_simple_sv_0_data_master_read),             //                                                .read
		.riscv_simple_sv_0_data_master_readdata                (riscv_simple_sv_0_data_master_readdata),         //                                                .readdata
		.riscv_simple_sv_0_data_master_readdatavalid           (riscv_simple_sv_0_data_master_readdatavalid),    //                                                .readdatavalid
		.riscv_simple_sv_0_data_master_write                   (riscv_simple_sv_0_data_master_write),            //                                                .write
		.riscv_simple_sv_0_data_master_writedata               (riscv_simple_sv_0_data_master_writedata),        //                                                .writedata
		.ledr_s1_address                                       (mm_interconnect_0_ledr_s1_address),              //                                         ledr_s1.address
		.ledr_s1_write                                         (mm_interconnect_0_ledr_s1_write),                //                                                .write
		.ledr_s1_readdata                                      (mm_interconnect_0_ledr_s1_readdata),             //                                                .readdata
		.ledr_s1_writedata                                     (mm_interconnect_0_ledr_s1_writedata),            //                                                .writedata
		.ledr_s1_chipselect                                    (mm_interconnect_0_ledr_s1_chipselect),           //                                                .chipselect
		.riscv_data_s1_address                                 (mm_interconnect_0_riscv_data_s1_address),        //                                   riscv_data_s1.address
		.riscv_data_s1_write                                   (mm_interconnect_0_riscv_data_s1_write),          //                                                .write
		.riscv_data_s1_readdata                                (mm_interconnect_0_riscv_data_s1_readdata),       //                                                .readdata
		.riscv_data_s1_writedata                               (mm_interconnect_0_riscv_data_s1_writedata),      //                                                .writedata
		.riscv_data_s1_byteenable                              (mm_interconnect_0_riscv_data_s1_byteenable),     //                                                .byteenable
		.riscv_data_s1_chipselect                              (mm_interconnect_0_riscv_data_s1_chipselect),     //                                                .chipselect
		.riscv_data_s1_clken                                   (mm_interconnect_0_riscv_data_s1_clken),          //                                                .clken
		.riscv_sdram_s1_address                                (mm_interconnect_0_riscv_sdram_s1_address),       //                                  riscv_sdram_s1.address
		.riscv_sdram_s1_write                                  (mm_interconnect_0_riscv_sdram_s1_write),         //                                                .write
		.riscv_sdram_s1_read                                   (mm_interconnect_0_riscv_sdram_s1_read),          //                                                .read
		.riscv_sdram_s1_readdata                               (mm_interconnect_0_riscv_sdram_s1_readdata),      //                                                .readdata
		.riscv_sdram_s1_writedata                              (mm_interconnect_0_riscv_sdram_s1_writedata),     //                                                .writedata
		.riscv_sdram_s1_byteenable                             (mm_interconnect_0_riscv_sdram_s1_byteenable),    //                                                .byteenable
		.riscv_sdram_s1_readdatavalid                          (mm_interconnect_0_riscv_sdram_s1_readdatavalid), //                                                .readdatavalid
		.riscv_sdram_s1_waitrequest                            (mm_interconnect_0_riscv_sdram_s1_waitrequest),   //                                                .waitrequest
		.riscv_sdram_s1_chipselect                             (mm_interconnect_0_riscv_sdram_s1_chipselect),    //                                                .chipselect
		.riscv_text_s1_address                                 (mm_interconnect_0_riscv_text_s1_address),        //                                   riscv_text_s1.address
		.riscv_text_s1_write                                   (mm_interconnect_0_riscv_text_s1_write),          //                                                .write
		.riscv_text_s1_readdata                                (mm_interconnect_0_riscv_text_s1_readdata),       //                                                .readdata
		.riscv_text_s1_writedata                               (mm_interconnect_0_riscv_text_s1_writedata),      //                                                .writedata
		.riscv_text_s1_byteenable                              (mm_interconnect_0_riscv_text_s1_byteenable),     //                                                .byteenable
		.riscv_text_s1_chipselect                              (mm_interconnect_0_riscv_text_s1_chipselect),     //                                                .chipselect
		.riscv_text_s1_clken                                   (mm_interconnect_0_riscv_text_s1_clken),          //                                                .clken
		.sw_s1_address                                         (mm_interconnect_0_sw_s1_address),                //                                           sw_s1.address
		.sw_s1_readdata                                        (mm_interconnect_0_sw_s1_readdata)                //                                                .readdata
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (sys_sdram_pll_reset_source_reset), // reset_in0.reset
		.clk            (sys_sdram_pll_sys_clk_clk),        //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),   // reset_out.reset
		.reset_req      (),                                 // (terminated)
		.reset_req_in0  (1'b0),                             // (terminated)
		.reset_in1      (1'b0),                             // (terminated)
		.reset_req_in1  (1'b0),                             // (terminated)
		.reset_in2      (1'b0),                             // (terminated)
		.reset_req_in2  (1'b0),                             // (terminated)
		.reset_in3      (1'b0),                             // (terminated)
		.reset_req_in3  (1'b0),                             // (terminated)
		.reset_in4      (1'b0),                             // (terminated)
		.reset_req_in4  (1'b0),                             // (terminated)
		.reset_in5      (1'b0),                             // (terminated)
		.reset_req_in5  (1'b0),                             // (terminated)
		.reset_in6      (1'b0),                             // (terminated)
		.reset_req_in6  (1'b0),                             // (terminated)
		.reset_in7      (1'b0),                             // (terminated)
		.reset_req_in7  (1'b0),                             // (terminated)
		.reset_in8      (1'b0),                             // (terminated)
		.reset_req_in8  (1'b0),                             // (terminated)
		.reset_in9      (1'b0),                             // (terminated)
		.reset_req_in9  (1'b0),                             // (terminated)
		.reset_in10     (1'b0),                             // (terminated)
		.reset_req_in10 (1'b0),                             // (terminated)
		.reset_in11     (1'b0),                             // (terminated)
		.reset_req_in11 (1'b0),                             // (terminated)
		.reset_in12     (1'b0),                             // (terminated)
		.reset_req_in12 (1'b0),                             // (terminated)
		.reset_in13     (1'b0),                             // (terminated)
		.reset_req_in13 (1'b0),                             // (terminated)
		.reset_in14     (1'b0),                             // (terminated)
		.reset_req_in14 (1'b0),                             // (terminated)
		.reset_in15     (1'b0),                             // (terminated)
		.reset_req_in15 (1'b0)                              // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (jtag_master_master_reset_reset),         // reset_in0.reset
		.reset_in1      (sys_sdram_pll_reset_source_reset),       // reset_in1.reset
		.clk            (sys_sdram_pll_sys_clk_clk),              //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_001_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

endmodule
